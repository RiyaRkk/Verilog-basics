module comparator(
  input [3:0]a,b,
  output out);
  assign out=(a>b);
endmodule
